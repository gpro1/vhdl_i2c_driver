%FDGF